library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL; 

entity processor is
  Port( clk: in STD_LOGIC;
        reset: in STD_LOGIC;
        start: in STD_LOGIC;
        
        Hready : in STD_LOGIC; --
        HRdata : in STD_LOGIC_VECTOR(31 downto 0); --
        
        Hwrite : out STD_LOGIC; --
        Haddr : out STD_LOGIC_VECTOR(15 downto 0); --
        Hsize : out STD_LOGIC_VECTOR(2 downto 0); --
        Htrans : out STD_LOGIC_VECTOR(1 downto 0); --
        HWdata : out STD_LOGIC_VECTOR(31 downto 0); --
        
        debug_controls : in STD_LOGIC_VECTOR(3 downto 0);
        debug_out : out STD_LOGIC_VECTOR(15 downto 0);
        ins_out : out STD_LOGIC_VECTOR(31 downto 0);
        Zout : out std_logic;
        Nout : out std_logic;
        Vout : out std_logic;
        Cout : out std_logic);
        --state : out STD_LOGIC_VECTOR(4 downto 0) );
end processor;

        
architecture Behavioral of processor is

    component controller
      Port(reset : in STD_LOGIC;
          clk : in STD_LOGIC;
          start : in STD_LOGIC;
          --control signals :
          carry : out STD_LOGIC;
          memoryReadEnable : out STD_LOGIC;
          memoryWriteEnable : out STD_LOGIC;
          IRenable : out STD_LOGIC;
          DRenable : out STD_LOGIC;
          RESenable : out STD_LOGIC;
          RFenable : out STD_LOGIC;
          Aenable : out STD_LOGIC;
          Benable : out STD_LOGIC;
          Menable : out STD_LOGIC;
          PMPathMode : out STD_LOGIC_VECTOR(2 downto 0);
          PMPathByteOffset : out STD_LOGIC_VECTOR(1 downto 0);
          ALUmode : out STD_LOGIC_VECTOR(3 downto 0);
          ALUop1select : out STD_LOGIC;
          ALUop2select : out STD_LOGIC_VECTOR(2 downto 0);
          rad1select : out STD_LOGIC_VECTOR(1 downto 0);
          rad2select : out STD_LOGIC;
          wadselect : out STD_LOGIC_VECTOR(1 downto 0);
          wdselect : out STD_LOGIC;
          Hwrite : out STD_LOGIC;
          Htrans : out STD_LOGIC_VECTOR(1 downto 0);
          --ShiftType : in STD_LOGIC_VECTOR(1 downto 0);  --read directly from instruction
          ShiftAmountSelect : out STD_LOGIC;
          ShifterInSelect : out STD_LOGIC;
          Fset : out STD_LOGIC;
          --output to controller :
          instruction : in STD_LOGIC_VECTOR(31 downto 0);
          Hready : in STD_LOGIC;
          flagZ : in STD_LOGIC;
          flagN : in STD_LOGIC;
          flagV : in STD_LOGIC;
          flagC : in STD_LOGIC;
          state_out : out STD_LOGIC_VECTOR(4 downto 0) );
    end component;
    
    component datapath
      Port (reset : in STD_LOGIC;
            clk : in STD_LOGIC;
            --control signals :
            carry : in STD_LOGIC;
            memoryReadEnable : in STD_LOGIC;
            memoryWriteEnable : in STD_LOGIC;
            IRenable : in STD_LOGIC;
            DRenable : in STD_LOGIC;
            RESenable : in STD_LOGIC;
            RFenable : in STD_LOGIC;
            Aenable : in STD_LOGIC;
            Benable : in STD_LOGIC;
            Menable : in STD_LOGIC;
            PMPathMode : in STD_LOGIC_VECTOR(2 downto 0);
            PMPathByteOffset : in STD_LOGIC_VECTOR(1 downto 0);
            ALUmode : in STD_LOGIC_VECTOR(3 downto 0);
            ALUop1select : in STD_LOGIC;
            ALUop2select : in STD_LOGIC_VECTOR(2 downto 0);
            rad1select : in STD_LOGIC_VECTOR(1 downto 0);
            rad2select : in STD_LOGIC;
            wadselect : in STD_LOGIC_VECTOR(1 downto 0);
            wdselect : in STD_LOGIC;
            HRdata : in STD_LOGIC_VECTOR(31 downto 0);
            --ShiftType : in STD_LOGIC_VECTOR(1 downto 0);  --read directly from instruction
            ShiftAmountSelect : in STD_LOGIC;
            ShifterInSelect : in STD_LOGIC;
            Fset : in STD_LOGIC;
            --output to controller :
            instruction : out STD_LOGIC_VECTOR(31 downto 0);
            flagZ : out STD_LOGIC;
            flagN : out STD_LOGIC;
            flagV : out STD_LOGIC;
            flagC : out STD_LOGIC;
            HWdata : out STD_LOGIC_VECTOR(31 downto 0);
            Haddr : out STD_LOGIC_VECTOR(15 downto 0);
            debug_controls : in STD_LOGIC_VECTOR(3 downto 0);
            debug_out : out STD_LOGIC_VECTOR(31 downto 0));
            
    end component;

    signal carry :  STD_LOGIC;
    signal memoryReadEnable :  STD_LOGIC;
    signal memoryWriteEnable :  STD_LOGIC;
    signal IRenable :  STD_LOGIC;
    signal DRenable :  STD_LOGIC;
    signal RESenable :  STD_LOGIC;
    signal RFenable :  STD_LOGIC;
    signal Aenable :  STD_LOGIC;
    signal Benable :  STD_LOGIC;
    signal Menable :  STD_LOGIC;
    signal PMPathMode :  STD_LOGIC_VECTOR(2 downto 0);
    signal PMPathByteOffset :  STD_LOGIC_VECTOR(1 downto 0);
    signal ALUmode :  STD_LOGIC_VECTOR(3 downto 0);
    signal ALUop1select :  STD_LOGIC;
    signal ALUop2select :  STD_LOGIC_VECTOR(2 downto 0);
    signal rad1select :  STD_LOGIC_VECTOR(1 downto 0);
    signal rad2select :  STD_LOGIC;
    signal wadselect :  STD_LOGIC_VECTOR(1 downto 0);
    signal wdselect :  STD_LOGIC;
    signal ShiftAmountSelect :  STD_LOGIC;
    signal ShifterSelect :  STD_LOGIC;
    signal Fset :  STD_LOGIC;
    signal instruction :  STD_LOGIC_VECTOR(31 downto 0);
    signal state_temp : STD_LOGIC_VECTOR(4 downto 0);
    signal flagZ :  STD_LOGIC;
    signal flagN :  STD_LOGIC;
    signal flagV :  STD_LOGIC;
    signal flagC :  STD_LOGIC;
    signal debug_out_internal : STD_LOGIC_VECTOR(31 downto 0) ;
begin

    Zout <= flagZ;
    Nout <= flagN;
    Vout <= flagV;
    Cout <= flagC;

    debug_out <= debug_out_internal(15 downto 0);
    ins_out <= instruction;
    
    Hsize <= "010";

    data_path: datapath
    Port Map(reset => reset,
            clk => clk,
            carry => carry,
            memoryReadEnable => memoryReadEnable,
            memoryWriteEnable => memoryWriteEnable,
            IRenable => IRenable,
            DRenable => DRenable,
            RESenable => RESenable,
            RFenable => RFenable,
            Aenable => Aenable,
            Benable => Benable,
            Menable => Menable,
            PMPathMode => PMPathMode,
            PMPathByteOffset => PMPathByteOffset,
            ALUmode => ALUmode,
            ALUop1select => ALUop1select,
            ALUop2select => ALUop2select,
            rad1select => rad1select,
            rad2select => rad2select,
            wadselect => wadselect,
            wdselect => wdselect,
            HRdata => HRdata,
            ShiftAmountSelect => ShiftAmountSelect,
            ShifterInSelect => ShifterSelect,
            Fset => Fset,
            instruction => instruction,
            flagZ => flagZ,
            flagN => flagN,
            flagV => flagV,
            flagC => flagC,
            HWdata => HWdata,
            Haddr => Haddr,
            debug_controls => debug_controls,
            debug_out => debug_out_internal);
            
    processor_controller: controller
    Port Map(reset => reset,
            clk => clk,
            start => start,
            carry => carry,
            memoryReadEnable => memoryReadEnable,
            memoryWriteEnable => memoryWriteEnable,
            IRenable => IRenable,
            DRenable => DRenable,
            RESenable => RESenable,
            RFenable => RFenable,
            Aenable => Aenable,
            Benable => Benable,
            Menable => Menable,
            PMPathMode => PMPathMode,
            PMPathByteOffset => PMPathByteOffset,
            ALUmode => ALUmode,
            ALUop1select => ALUop1select,
            ALUop2select => ALUop2select,
            rad1select => rad1select,
            rad2select => rad2select,
            wadselect => wadselect,
            wdselect => wdselect,
            Hwrite => Hwrite,
            Htrans => Htrans,
            ShiftAmountSelect => ShiftAmountSelect,
            ShifterInSelect => ShifterSelect,
            Fset => Fset,
            instruction => instruction,
            Hready => Hready,
            flagZ => flagZ,
            flagN => flagN,
            flagV => flagV,
            flagC => flagC,
            state_out => state_temp);
            
    --state <= state_temp;

end architecture;